library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

entity function_R is
    generic ( N : INTEGER := 41);
    port (
        input_vector            : in std_logic_vector (N - 1 downto 0);
        output_result : out std_logic_vector(N+N-2 downto 0)
        );
end function_R;
architecture behavorial of function_R is
begin
    process(input_vector)
    begin
        if input_vector(0) = '1' then
            output_result(0) <= '1';
        else
            output_result(0) <= '0';
        end if;

        if input_vector(1) = '1' then
            output_result(1) <= '1';
        else
            output_result(1) <= '0';
        end if;

        if input_vector(2) = '1' then
            output_result(2) <= '1';
        else
            output_result(2) <= '0';
        end if;

        if input_vector(3) = '1' then
            output_result(3) <= '1';
        else
            output_result(3) <= '0';
        end if;

        if input_vector(4) = '1' then
            output_result(4) <= '1';
        else
            output_result(4) <= '0';
        end if;

        if input_vector(5) = '1' then
            output_result(5) <= '1';
        else
            output_result(5) <= '0';
        end if;

        if input_vector(6) = '1' then
            output_result(6) <= '1';
        else
            output_result(6) <= '0';
        end if;

        if input_vector(7) = '1' then
            output_result(7) <= '1';
        else
            output_result(7) <= '0';
        end if;

        if input_vector(8) = '1' then
            output_result(8) <= '1';
        else
            output_result(8) <= '0';
        end if;

        if input_vector(9) = '1' then
            output_result(9) <= '1';
        else
            output_result(9) <= '0';
        end if;

        if input_vector(10) = '1' then
            output_result(10) <= '1';
        else
            output_result(10) <= '0';
        end if;

        if input_vector(11) = '1' then
            output_result(11) <= '1';
        else
            output_result(11) <= '0';
        end if;

        if input_vector(11) = '1' then
            output_result(11) <= '1';
        else
            output_result(11) <= '0';
        end if;

        if input_vector(12) = '1' then
            output_result(12) <= '1';
        else
            output_result(12) <= '0';
        end if;

        if input_vector(13) = '1' then
            output_result(13) <= '1';
        else
            output_result(13) <= '0';
        end if;

        if input_vector(14) = '1' then
            output_result(14) <= '1';
        else
            output_result(14) <= '0';
        end if;

        if input_vector(15) = '1' then
            output_result(15) <= '1';
        else
            output_result(15) <= '0';
        end if;

        if input_vector(16) = '1' then
            output_result(16) <= '1';
        else
            output_result(16) <= '0';
        end if;

        if input_vector(17) = '1' then
            output_result(17) <= '1';
        else
            output_result(17) <= '0';
        end if;

        if input_vector(18) = '1' then
            output_result(18) <= '1';
        else
            output_result(18) <= '0';
        end if;

        if input_vector(19) = '1' then
            output_result(19) <= '1';
        else
            output_result(19) <= '0';
        end if;

        if input_vector(20) = '1' then
            output_result(20) <= '1';
        else
            output_result(20) <= '0';
        end if;

        if input_vector(21) = '1' then
            output_result(21) <= '1';
        else
            output_result(21) <= '0';
        end if;

        if input_vector(22) = '1' then
            output_result(22) <= '1';
        else
            output_result(22) <= '0';
        end if;

        if input_vector(23) = '1' then
            output_result(23) <= '1';
        else
            output_result(23) <= '0';
        end if;

        if input_vector(24) = '1' then
            output_result(24) <= '1';
        else
            output_result(24) <= '0';
        end if;

        if input_vector(25) = '1' then
            output_result(25) <= '1';
        else
            output_result(25) <= '0';
        end if;

        if input_vector(26) = '1' then
            output_result(26) <= '1';
        else
            output_result(26) <= '0';
        end if;

        if input_vector(27) = '1' then
            output_result(27) <= '1';
        else
            output_result(27) <= '0';
        end if;

        if input_vector(28) = '1' then
            output_result(28) <= '1';
        else
            output_result(28) <= '0';
        end if;

        if input_vector(29) = '1' then
            output_result(29) <= '1';
        else
            output_result(29) <= '0';
        end if;

        if input_vector(30) = '1' then
            output_result(30) <= '1';
        else
            output_result(30) <= '0';
        end if;

        if input_vector(31) = '1' then
            output_result(31) <= '1';
        else
            output_result(31) <= '0';
        end if;

        if input_vector(32) = '1' then
            output_result(32) <= '1';
        else
            output_result(32) <= '0';
        end if;

        if input_vector(33) = '1' then
            output_result(33) <= '1';
        else
            output_result(33) <= '0';
        end if;

        if input_vector(34) = '1' then
            output_result(34) <= '1';
        else
            output_result(34) <= '0';
        end if;

        if input_vector(35) = '1' then
            output_result(35) <= '1';
        else
            output_result(35) <= '0';
        end if;

        if input_vector(36) = '1' then
            output_result(36) <= '1';
        else
            output_result(36) <= '0';
        end if;

        if input_vector(37) = '1' then
            output_result(37) <= '1';
        else
            output_result(37) <= '0';
        end if;

        
        if input_vector(38) = '1' then
            output_result(38) <= '1';
        else
            output_result(38) <= '0';
        end if;

        
        if input_vector(39) = '1' then
            output_result(39) <= '1';
        else
            output_result(39) <= '0';
        end if;

        output_result(80 downto 40) <= (others => '0');
    end process;
end behavorial;

