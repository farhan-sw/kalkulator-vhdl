library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity KalkulatorTopLevel is
	generic ( N : Integer := 41);
	port (
		P, Q		: IN STD_LOGIC_VECTOR (N-1 DOWNTO 0);
		M 			: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		CLK 		: IN STD_LOGIC;
		RST			: IN STD_LOGIC;
		OUT_OPERASI	: OUT STD_LOGIC_VECTOR (N-1 DOWNTO 0);
		STATUS 		: OUT STD_LOGIC_VECTOR (1 DOWNTO 0)
	);
end KalkulatorTopLevel;


architecture KalkulatorTopLevel_arc of KalkulatorTopLevel is 

component AdderSubtractor is
    generic ( N : INTEGER := N);
    port (
        P_in            : in std_logic_vector (N - 1 downto 0);
        Q_in            : in std_logic_vector (N - 1 downto 0);

        OUT_Operasi     : out std_logic_vector (N - 1 downto 0);

        M               : in std_logic_vector(2 downto 0);
        status          : out std_logic_vector(1 downto 0);

        clk             : in std_logic;
        rst             : in std_logic
    );
end component;


component divider is
    generic ( N : INTEGER := N);
    port (
        P_in            : in std_logic_vector (N - 1 downto 0);
        Q_in            : in std_logic_vector (N - 1 downto 0);

        ---OUT_Operasi     : buffer std_logic_vector (N - 1 downto 0);
        out_operasi_fix : out std_logic_vector (N - 1 downto 0);

        M               : in std_logic_vector(2 downto 0);
        status          : out std_logic_vector(1 downto 0);

		debug_fsm : out std_logic_vector(3 downto 0);
		debug_m1, debug_m2 : out std_logic_vector (N-1 downto 0);
        clk             : in std_logic;
        rst             : in std_logic
    );
end component;

component FPB is 
	generic ( N: INTEGER := N);
	port (
		P_in, Q_in : IN STD_LOGIC_VECTOR (N-1 downto 0);
		Mode : IN STD_LOGIC_VECTOR (2 downto 0);
		St : OUT STD_LOGIC_VECTOR (1 downto 0); 
		OUT_FPB: OUT STD_LOGIC_VECTOR (N-1 downto 0); 
        clk, rst : IN STD_LOGIC );
end component;


component Multiplication is 
	generic ( N: INTEGER := N);
	port (
		P			: in std_logic_vector (N-1 downto 0) ;
		Q			: in std_logic_vector (N-1 downto 0) ;
		Mode		: in std_logic_vector (2 downto 0) ;
		Clk, Rst	: in std_logic ;
		Multi_Out	: out std_logic_vector (N-1 downto 0) ;
		Status_Out	: out std_logic_vector (1 downto 0) ;
		debugout 	: out integer 
	);
end component;

component Pangkat is  
	generic ( N: INTEGER := 41); 
	port ( 
		P_in   	      : in std_logic_vector (N-1 downto 0); 
		Q_in          : in std_logic_vector (N-1 downto 0); 
		Mode          : in std_logic_vector (2 downto 0); 

        clk           : in std_logic; 
        rst           : in std_logic; 

		out_pangkat   : out std_logic_vector (N-1 downto 0);  
		status        : out std_logic_vector (1 downto 0);  

        debug_pangkat : out integer
	); 
end component; 


component mux8to1 is
    generic ( N : INTEGER := N);
    port (
        IN1                  : in std_logic_vector (N-1 downto 0);
        IN2                  : in std_logic_vector (N-1 downto 0);
        IN3                  : in std_logic_vector (N-1 downto 0);
        IN4                  : in std_logic_vector (N-1 downto 0);
        IN5                  : in std_logic_vector (N-1 downto 0);
        IN6                  : in std_logic_vector (N-1 downto 0);
        IN7                  : in std_logic_vector (N-1 downto 0);

        S                    : in std_logic_vector (2 downto 0);
        OUTMUX               : out std_logic_vector(N-1 downto 0);

        clk                  : in std_logic

    );
end component;

component mux8to1stat is
    port (
        IN1                  : in std_logic_vector (1 downto 0);
        IN2                  : in std_logic_vector (1 downto 0);
        IN3                  : in std_logic_vector (1 downto 0);
        IN4                  : in std_logic_vector (1 downto 0);
        IN5                  : in std_logic_vector (1 downto 0);
        IN6                  : in std_logic_vector (1 downto 0);
        IN7                  : in std_logic_vector (1 downto 0);

        S                    : in std_logic_vector (2 downto 0);
        OUTMUX               : out std_logic_vector(1 downto 0);

        clk                  : in std_logic

    );
end component;

signal outAdderSubtractor, outdivider, outFPB, outOperasi, outMulti, outPangkat  : std_logic_vector (N-1 downto 0);
signal statAdderSubtractor, statdivider, statFPB, statOutput, statMulti, statPangkat : std_logic_vector (1 downto 0);
signal kosongkeluar : std_logic_vector (N-1 downto 0) := (others => '0');
signal kosongstatus : std_logic_vector (1 downto 0) := "00";
signal debug_fsmm : std_logic_vector (3 downto 0); 
signal debug_m11, debug_m22 : std_logic_vector (N-1 downto 0);
signal debugg,debugs : integer;

begin

	blockAdderSubtractor : AdderSubtractor port map (P, Q, outAdderSubtractor, M, statAdderSubtractor, clk, rst);
	blockdivider : divider port map (P, Q, outdivider, M, statdivider, debug_fsmm, debug_m11, debug_m22, clk, rst);
	blockFPB : FPB port map (P, Q, M, statFPB, outFPB, clk, rst);
	blockMulti : multiplication port map (P, Q, M, clk, rst, outMulti, statmulti, debugg);
	blockPangkat : Pangkat port map (P, Q, M, clk ,rst, outPangkat, statPangkat, debugs);
	
	mux8to1Out : mux8to1 port map (outAdderSubtractor,outAdderSubtractor,outMulti, outdivider, outdivider, outPangkat, outFPB,  M, outOperasi, clk);
	mux8to1Stats : mux8to1stat port map ( statAdderSubtractor, statAdderSubtractor, statMulti, statdivider, statdivider, statPangkat, statFPB, M, statOutput, clk);
	
	process (clk)
	begin
		OUT_Operasi <= outOperasi;
		status <= statOutput;
	end process; 
	
end KalkulatorTopLevel_arc;

